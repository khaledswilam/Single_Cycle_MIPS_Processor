module sh_left32(input [31:0] in32,
output [31:0] out32);
 
     
   
	   
      assign out32=in32<<2;

     
	
 
endmodule